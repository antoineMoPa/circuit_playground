* sim.spice

.get circuit.net

.print op v(4) i(RL)

.op
